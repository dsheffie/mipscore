module fpu (
	clk,
	reset,
	pc,
	opcode,
	start,
	src_a,
	src_b,
	src_c,
	src_fcr,
	rob_ptr_in,
	dst_ptr_in,
	fcr_ptr_in,
	fcr_sel,
	val,
	cmp_val,
	y,
	rob_ptr_out,
	dst_ptr_out,
	fcr_ptr_out
);
	parameter LG_PRF_WIDTH = 4;
	parameter LG_ROB_WIDTH = 4;
	parameter LG_FCR_WIDTH = 4;
	parameter FPU_LAT = 2;
	input wire clk;
	input wire reset;
	input wire [63:0] pc;
	input opcode_t opcode;
	input wire start;
	input wire [63:0] src_a;
	input wire [63:0] src_b;
	input wire [63:0] src_c;
	input wire [7:0] src_fcr;
	input wire [LG_ROB_WIDTH - 1:0] rob_ptr_in;
	input wire [LG_PRF_WIDTH - 1:0] dst_ptr_in;
	input wire [LG_FCR_WIDTH - 1:0] fcr_ptr_in;
	input wire [2:0] fcr_sel;
	output reg val;
	output reg cmp_val;
	output reg [63:0] y;
	output wire [LG_ROB_WIDTH - 1:0] rob_ptr_out;
	output wire [LG_PRF_WIDTH - 1:0] dst_ptr_out;
	output wire [LG_FCR_WIDTH - 1:0] fcr_ptr_out;
	wire [31:0] t_sp_adder_result;
	wire [63:0] t_dp_adder_result;
	wire [31:0] t_sp_mult_result;
	wire [63:0] t_dp_mult_result;
	reg [FPU_LAT - 1:0] r_val;
	reg [LG_PRF_WIDTH - 1:0] r_ptr [FPU_LAT - 1:0];
	reg [LG_ROB_WIDTH - 1:0] r_rob [FPU_LAT - 1:0];
	reg [LG_FCR_WIDTH - 1:0] r_fcr [FPU_LAT - 1:0];
	reg [2:0] r_fcr_sel [FPU_LAT - 1:0];
	reg [7:0] r_fcr_reg [FPU_LAT - 1:0];
	wire [7:0] fcr_reg;
	opcode_t r_opcode [FPU_LAT - 1:0];
	assign dst_ptr_out = r_ptr[0];
	assign rob_ptr_out = r_rob[0];
	assign fcr_ptr_out = r_fcr[0];
	assign fcr_reg = r_fcr_reg[0];
	wire w_sp_cmp;
	wire w_dp_cmp;
	reg [3:0] t_sp_cmp_type;
	reg [3:0] t_dp_cmp_type;
	always @(*) begin
		t_sp_cmp_type = 4'd0;
		case (opcode)
			SP_CMP_LT: t_sp_cmp_type = 4'd1;
			SP_CMP_EQ: t_sp_cmp_type = 4'd3;
			SP_CMP_LE: t_sp_cmp_type = 4'd2;
			default:
				;
		endcase
	end
	always @(*) begin
		t_dp_cmp_type = 4'd0;
		case (opcode)
			DP_CMP_LT: t_dp_cmp_type = 4'd1;
			DP_CMP_EQ: t_dp_cmp_type = 4'd3;
			DP_CMP_LE: t_dp_cmp_type = 4'd2;
			default:
				;
		endcase
	end
	fp_compare #(
		.W(32),
		.D(FPU_LAT)
	) sp_cmp(
		.clk(clk),
		.pc(pc),
		.a(src_a[31:0]),
		.b(src_b[31:0]),
		.start(start && (t_sp_cmp_type != 4'd0)),
		.cmp_type(t_sp_cmp_type),
		.y(w_sp_cmp)
	);
	fp_compare #(
		.W(64),
		.D(FPU_LAT)
	) dp_cmp(
		.clk(clk),
		.pc(pc),
		.a(src_a),
		.b(src_b),
		.start(start && (t_dp_cmp_type != 4'd0)),
		.cmp_type(t_dp_cmp_type),
		.y(w_dp_cmp)
	);
	function [63:0] handle_fcr;
		input reg b;
		input reg [2:0] sel;
		input reg [7:0] fcr_reg;
		reg [63:0] y;
		begin
			case (sel)
				3'd0: y = {56'd0, fcr_reg[7:1], b};
				3'd1: y = {56'd0, fcr_reg[7:2], b, fcr_reg[0]};
				3'd2: y = {56'd0, fcr_reg[7:3], b, fcr_reg[1:0]};
				3'd3: y = {56'd0, fcr_reg[7:4], b, fcr_reg[2:0]};
				3'd4: y = {56'd0, fcr_reg[7:5], b, fcr_reg[3:0]};
				3'd5: y = {56'd0, fcr_reg[7:6], b, fcr_reg[4:0]};
				3'd6: y = {56'd0, fcr_reg[7], b, fcr_reg[5:0]};
				3'd7: y = {56'd0, b, fcr_reg[6:0]};
			endcase
			handle_fcr = y;
		end
	endfunction
	always @(*) begin
		y = 'd0;
		val = 1'b0;
		cmp_val = 1'b0;
		case (r_opcode[0])
			SP_ADD: begin
				y = {32'd0, t_sp_adder_result};
				val = r_val[0];
			end
			SP_SUB: begin
				y = {32'd0, t_sp_adder_result};
				val = r_val[0];
			end
			DP_ADD: begin
				y = t_dp_adder_result;
				val = r_val[0];
			end
			DP_SUB: begin
				y = t_dp_adder_result;
				val = r_val[0];
			end
			SP_MUL: begin
				y = {32'd0, t_sp_mult_result};
				val = r_val[0];
			end
			DP_MUL: begin
				y = t_dp_mult_result;
				val = r_val[0];
			end
			SP_CMP_LT: begin
				cmp_val = r_val[0];
				y = handle_fcr(w_sp_cmp, r_fcr_sel[0], fcr_reg);
			end
			SP_CMP_LE: begin
				cmp_val = r_val[0];
				y = handle_fcr(w_sp_cmp, r_fcr_sel[0], fcr_reg);
			end
			SP_CMP_EQ: begin
				cmp_val = r_val[0];
				y = handle_fcr(w_sp_cmp, r_fcr_sel[0], fcr_reg);
			end
			DP_CMP_LT: begin
				cmp_val = r_val[0];
				y = handle_fcr(w_dp_cmp, r_fcr_sel[0], fcr_reg);
			end
			DP_CMP_LE: begin
				cmp_val = r_val[0];
				y = handle_fcr(w_dp_cmp, r_fcr_sel[0], fcr_reg);
			end
			DP_CMP_EQ: begin
				cmp_val = r_val[0];
				y = handle_fcr(w_dp_cmp, r_fcr_sel[0], fcr_reg);
			end
			default:
				;
		endcase
	end
	always @(posedge clk)
		if (reset)
			r_val <= 'd0;
		else begin
			r_val[FPU_LAT - 1] <= start;
			begin : sv2v_autoblock_1
				integer i;
				for (i = FPU_LAT - 1; i > 0; i = i - 1)
					r_val[i - 1] <= r_val[i];
			end
		end
	always @(posedge clk) begin
		r_opcode[FPU_LAT - 1] <= opcode;
		r_ptr[FPU_LAT - 1] <= dst_ptr_in;
		r_fcr[FPU_LAT - 1] <= fcr_ptr_in;
		r_rob[FPU_LAT - 1] <= rob_ptr_in;
		r_fcr_sel[FPU_LAT - 1] <= fcr_sel;
		r_fcr_reg[FPU_LAT - 1] <= src_fcr;
		begin : sv2v_autoblock_2
			integer i;
			for (i = FPU_LAT - 1; i > 0; i = i - 1)
				begin
					r_opcode[i - 1] <= r_opcode[i];
					r_ptr[i - 1] <= r_ptr[i];
					r_fcr[i - 1] <= r_fcr[i];
					r_rob[i - 1] <= r_rob[i];
					r_fcr_sel[i - 1] <= r_fcr_sel[i];
					r_fcr_reg[i - 1] <= r_fcr_reg[i];
				end
		end
	end
	fp_add #(
		.W(32),
		.ADD_LAT(FPU_LAT)
	) sa(
		.clk(clk),
		.sub(opcode == SP_SUB),
		.a(src_a[31:0]),
		.b(src_b[31:0]),
		.en((opcode == SP_ADD) || (opcode == SP_SUB)),
		.y(t_sp_adder_result)
	);
	fp_add #(
		.W(64),
		.ADD_LAT(FPU_LAT)
	) sd(
		.clk(clk),
		.sub(opcode == DP_SUB),
		.a(src_a),
		.b(src_b),
		.en((opcode == DP_ADD) || (opcode == DP_SUB)),
		.y(t_dp_adder_result)
	);
	fp_mul #(
		.W(32),
		.MUL_LAT(FPU_LAT)
	) sm(
		.clk(clk),
		.a(src_a[31:0]),
		.b(src_b[31:0]),
		.en(opcode == SP_MUL),
		.y(t_sp_mult_result)
	);
	fp_mul #(
		.W(64),
		.MUL_LAT(FPU_LAT)
	) dm(
		.clk(clk),
		.a(src_a[63:0]),
		.b(src_b[63:0]),
		.en(opcode == DP_MUL),
		.y(t_dp_mult_result)
	);
endmodule
